module unidade_logica(
	input [2:0] operacao,
	input [224:0] matriz_A,
	input [224:0] matriz_B,
	output reg [224:0] matriz_resultado,
);
	
	
			
endmodule